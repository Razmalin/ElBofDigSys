rom_1_inst : rom_1 PORT MAP (
		address	 => address_sig,
		inclock	 => inclock_sig,
		outclock	 => outclock_sig,
		q	 => q_sig
	);
